* AD820  SPICE Macro-model                 
* Description: Amplifier
* Generic Desc: 5/30V, JFET, OP, S SPLY, RRO, 1X
* Developed by: JCB / PMI
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (08/1991)
* Copyright 1993, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node assignments
*                non-inverting input
*                | inverting input
*                | | positive supply
*                | | |  negative supply
*                | | |  |  output
*                | | |  |  |
.SUBCKT AD820    1 2 99 50 25
*
* INPUT STAGE & POLE AT 3 MHZ
*
R3   5  99   2456
R4   6  99   2456
CIN  1   2   5E-12
C2   5   6   10.8E-12
I1   4  50   108E-6
IOS  1   2   1E-12
EOS  7   1   POLY(1) (12,98) 100E-6  1
J1   4   2   5   JX
J2   4   7   6   JX
*
EREF 98  0   30  0  1
*
* GAIN STAGE & POLE AT 124 HZ
*
R5   9  98   2.46E6
C3   9  25   35E-12
G1   98  9   6  5  4.07E-4
V1   8  98   0
V2   98 10   -1
D1   9  10   DX
D2   8   9   DX
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 1 KHZ
*
R21  11 12   1E6
R22  12 98   1
C14  11 12   159E-12
E13  11 98   POLY(2) (2,98) (1,98) 0 50 50
*
* POLE AT 10 MHZ
*
R23  18 98   1E6
C15  18 98   15.9E-15
G15  98 18   9  98  1E-6
*
* OUTPUT STAGE
*
ES   26  51  POLY(1) (18,98) 1.72 1
RS   26  22  500
V3   23  51  1.1
V4   21  23  1.36
C16  20  25  2E-12
C17  24  25  2E-12
RG1  20  97  1E8
RG2  24  97  1E8
Q1   20  20  97  PNP
Q2   20  21  22  NPN
Q3   24  23  22  PNP
Q4   24  24  51  NPN
Q5   25  20  97  PNP 20
Q6   25  24  51  NPN 20
VP   96  97  0
VN   51  52  0
EP   96  0   POLY(1) (99,0) 0.01 1
EN   52  0   POLY(1) (50,0) -0.015 1
*
R25  30 99   5E6
R26  30 50   5E6
FSY1 99  0   VP 1
FSY2 0  50   VN 1 
*
* MODELS USED
*
.MODEL JX   NJF(BETA=7.67E-4  VTO=-2.000  IS=1E-12)
.MODEL NPN  NPN(BF=120 VAF=150 VAR=15 RB=2E3
+ RE=4 RC=200 IS=1E-16)
.MODEL PNP  PNP(BF=80 VAF=150 VAR=15 RB=2E3
+ RE=4 RC=900 IS=1E-16)
.MODEL DX   D(IS=1E-15)
.ENDS AD820





